// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// Generated by Quartus Prime Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition
// Created on Tue Nov 16 18:53:44 2021

// synthesis message_off 10175

`timescale 1ns/1ns

module test (
    reset,clock,Din,
    correct);

    input reset;
    input clock;
    input [3:0] Din;
    tri0 reset;
    tri0 [3:0] Din;
    output correct;
    reg correct;
    reg [4:0] fstate;
    reg [4:0] reg_fstate;
    parameter state1=0,state2=1,state3=2,state4=3,state5=4;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or Din)
    begin
        if (~reset) begin
            reg_fstate <= state1;
            correct <= 1'b0;
        end
        else begin
            correct <= 1'b0;
            case (fstate)
                state1: begin
                    if ((Din[3:0] != 4'b0100))
                        reg_fstate <= state1;
                    else if ((Din[3:0] == 4'b0100))
                        reg_fstate <= state2;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state1;

                    correct <= 1'b0;
                end
                state2: begin
                    if ((Din[3:0] != 4'b0101))
                        reg_fstate <= state1;
                    else if ((Din[3:0] == 4'b0101))
                        reg_fstate <= state3;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state2;

                    correct <= 1'b0;
                end
                state3: begin
                    if ((Din[3:0] != 4'b0111))
                        reg_fstate <= state1;
                    else if ((Din[3:0] == 4'b0111))
                        reg_fstate <= state4;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state3;

                    correct <= 1'b0;
                end
                state4: begin
                    if ((Din[3:0] != 4'b1001))
                        reg_fstate <= state1;
                    else if ((Din[3:0] == 4'b1001))
                        reg_fstate <= state5;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state4;

                    correct <= 1'b0;
                end
                state5: begin
                    if ((Din[3:0] != 4'b0100))
                        reg_fstate <= state1;
                    else if ((Din[3:0] == 4'b0100))
                        reg_fstate <= state2;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state5;

                    correct <= 1'b1;
                end
                default: begin
                    correct <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // test
