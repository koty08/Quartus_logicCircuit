// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition"
// CREATED		"Wed Dec 22 12:35:05 2021"

module ascii_comparator(
	ASCII_Input,
	is_ADD,
	is_SUB,
	is_MOV,
	is_SHW
);


input wire	[7:0] ASCII_Input;
output wire	is_ADD;
output wire	is_SUB;
output wire	is_MOV;
output wire	is_SHW;

wire	[7:0] l_input;
wire	SYNTHESIZED_WIRE_0;
wire	SYNTHESIZED_WIRE_1;
wire	SYNTHESIZED_WIRE_2;
wire	SYNTHESIZED_WIRE_3;
wire	SYNTHESIZED_WIRE_4;
wire	SYNTHESIZED_WIRE_5;
wire	SYNTHESIZED_WIRE_6;
wire	SYNTHESIZED_WIRE_7;
wire	SYNTHESIZED_WIRE_8;
wire	SYNTHESIZED_WIRE_9;
wire	SYNTHESIZED_WIRE_10;
wire	SYNTHESIZED_WIRE_11;
wire	SYNTHESIZED_WIRE_12;
wire	SYNTHESIZED_WIRE_91;
wire	SYNTHESIZED_WIRE_20;
wire	SYNTHESIZED_WIRE_22;
wire	SYNTHESIZED_WIRE_24;
wire	SYNTHESIZED_WIRE_26;
wire	SYNTHESIZED_WIRE_27;
wire	SYNTHESIZED_WIRE_28;
wire	SYNTHESIZED_WIRE_29;
wire	SYNTHESIZED_WIRE_30;
wire	SYNTHESIZED_WIRE_31;
wire	SYNTHESIZED_WIRE_32;
wire	SYNTHESIZED_WIRE_33;
wire	SYNTHESIZED_WIRE_34;
wire	SYNTHESIZED_WIRE_35;
wire	SYNTHESIZED_WIRE_40;
wire	SYNTHESIZED_WIRE_42;
wire	SYNTHESIZED_WIRE_43;
wire	SYNTHESIZED_WIRE_44;
wire	SYNTHESIZED_WIRE_49;
wire	SYNTHESIZED_WIRE_50;
wire	SYNTHESIZED_WIRE_51;
wire	SYNTHESIZED_WIRE_52;
wire	SYNTHESIZED_WIRE_53;
wire	SYNTHESIZED_WIRE_54;
wire	SYNTHESIZED_WIRE_55;
wire	SYNTHESIZED_WIRE_56;
wire	SYNTHESIZED_WIRE_57;
wire	SYNTHESIZED_WIRE_58;
wire	SYNTHESIZED_WIRE_63;
wire	SYNTHESIZED_WIRE_65;
wire	SYNTHESIZED_WIRE_66;
wire	SYNTHESIZED_WIRE_68;
wire	SYNTHESIZED_WIRE_69;
wire	SYNTHESIZED_WIRE_70;
wire	SYNTHESIZED_WIRE_71;
wire	SYNTHESIZED_WIRE_72;
wire	SYNTHESIZED_WIRE_73;
wire	SYNTHESIZED_WIRE_74;
wire	SYNTHESIZED_WIRE_75;
wire	SYNTHESIZED_WIRE_76;
wire	SYNTHESIZED_WIRE_77;
wire	SYNTHESIZED_WIRE_78;
wire	SYNTHESIZED_WIRE_79;
wire	SYNTHESIZED_WIRE_80;
wire	SYNTHESIZED_WIRE_81;
wire	SYNTHESIZED_WIRE_88;
wire	SYNTHESIZED_WIRE_89;

assign	SYNTHESIZED_WIRE_91 = 1;




assign	SYNTHESIZED_WIRE_9 = l_input[1] ~^ SYNTHESIZED_WIRE_0;

assign	SYNTHESIZED_WIRE_10 = l_input[0] ~^ SYNTHESIZED_WIRE_1;

assign	SYNTHESIZED_WIRE_26 = l_input[7] ~^ SYNTHESIZED_WIRE_2;

assign	SYNTHESIZED_WIRE_11 = SYNTHESIZED_WIRE_3 & SYNTHESIZED_WIRE_4 & SYNTHESIZED_WIRE_5 & SYNTHESIZED_WIRE_6;

assign	SYNTHESIZED_WIRE_12 = SYNTHESIZED_WIRE_7 & SYNTHESIZED_WIRE_8 & SYNTHESIZED_WIRE_9 & SYNTHESIZED_WIRE_10;

assign	is_ADD = SYNTHESIZED_WIRE_11 & SYNTHESIZED_WIRE_12;

assign	SYNTHESIZED_WIRE_44 =  ~SYNTHESIZED_WIRE_91;

assign	SYNTHESIZED_WIRE_79 =  ~SYNTHESIZED_WIRE_91;

assign	SYNTHESIZED_WIRE_88 =  ~SYNTHESIZED_WIRE_91;

assign	SYNTHESIZED_WIRE_89 =  ~SYNTHESIZED_WIRE_91;

assign	SYNTHESIZED_WIRE_0 =  ~SYNTHESIZED_WIRE_91;

assign	SYNTHESIZED_WIRE_1 =  ~SYNTHESIZED_WIRE_91;

assign	SYNTHESIZED_WIRE_27 = l_input[6] ~^ SYNTHESIZED_WIRE_91;

assign	SYNTHESIZED_WIRE_28 = l_input[5] ~^ SYNTHESIZED_WIRE_20;

assign	SYNTHESIZED_WIRE_29 = l_input[4] ~^ SYNTHESIZED_WIRE_91;

assign	SYNTHESIZED_WIRE_30 = l_input[3] ~^ SYNTHESIZED_WIRE_22;

assign	SYNTHESIZED_WIRE_31 = l_input[2] ~^ SYNTHESIZED_WIRE_91;

assign	SYNTHESIZED_WIRE_32 = l_input[1] ~^ SYNTHESIZED_WIRE_24;

assign	SYNTHESIZED_WIRE_33 = l_input[0] ~^ SYNTHESIZED_WIRE_91;

assign	SYNTHESIZED_WIRE_34 = SYNTHESIZED_WIRE_26 & SYNTHESIZED_WIRE_27 & SYNTHESIZED_WIRE_28 & SYNTHESIZED_WIRE_29;

assign	SYNTHESIZED_WIRE_35 = SYNTHESIZED_WIRE_30 & SYNTHESIZED_WIRE_31 & SYNTHESIZED_WIRE_32 & SYNTHESIZED_WIRE_33;

assign	is_SUB = SYNTHESIZED_WIRE_34 & SYNTHESIZED_WIRE_35;

assign	SYNTHESIZED_WIRE_2 =  ~SYNTHESIZED_WIRE_91;

assign	SYNTHESIZED_WIRE_20 =  ~SYNTHESIZED_WIRE_91;

assign	SYNTHESIZED_WIRE_22 =  ~SYNTHESIZED_WIRE_91;

assign	SYNTHESIZED_WIRE_24 =  ~SYNTHESIZED_WIRE_91;

assign	SYNTHESIZED_WIRE_49 = l_input[7] ~^ SYNTHESIZED_WIRE_40;

assign	SYNTHESIZED_WIRE_50 = l_input[6] ~^ SYNTHESIZED_WIRE_91;

assign	SYNTHESIZED_WIRE_51 = l_input[5] ~^ SYNTHESIZED_WIRE_42;

assign	SYNTHESIZED_WIRE_52 = l_input[4] ~^ SYNTHESIZED_WIRE_43;

assign	SYNTHESIZED_WIRE_3 = l_input[7] ~^ SYNTHESIZED_WIRE_44;

assign	SYNTHESIZED_WIRE_53 = l_input[3] ~^ SYNTHESIZED_WIRE_91;

assign	SYNTHESIZED_WIRE_54 = l_input[2] ~^ SYNTHESIZED_WIRE_91;

assign	SYNTHESIZED_WIRE_55 = l_input[1] ~^ SYNTHESIZED_WIRE_91;

assign	SYNTHESIZED_WIRE_56 = l_input[0] ~^ SYNTHESIZED_WIRE_91;

assign	SYNTHESIZED_WIRE_57 = SYNTHESIZED_WIRE_49 & SYNTHESIZED_WIRE_50 & SYNTHESIZED_WIRE_51 & SYNTHESIZED_WIRE_52;

assign	SYNTHESIZED_WIRE_58 = SYNTHESIZED_WIRE_53 & SYNTHESIZED_WIRE_54 & SYNTHESIZED_WIRE_55 & SYNTHESIZED_WIRE_56;

assign	is_MOV = SYNTHESIZED_WIRE_57 & SYNTHESIZED_WIRE_58;

assign	SYNTHESIZED_WIRE_40 =  ~SYNTHESIZED_WIRE_91;

assign	SYNTHESIZED_WIRE_42 =  ~SYNTHESIZED_WIRE_91;

assign	SYNTHESIZED_WIRE_43 =  ~SYNTHESIZED_WIRE_91;

assign	SYNTHESIZED_WIRE_4 = l_input[6] ~^ SYNTHESIZED_WIRE_91;

assign	SYNTHESIZED_WIRE_71 = l_input[7] ~^ SYNTHESIZED_WIRE_63;

assign	SYNTHESIZED_WIRE_72 = l_input[6] ~^ SYNTHESIZED_WIRE_91;

assign	SYNTHESIZED_WIRE_73 = l_input[5] ~^ SYNTHESIZED_WIRE_65;

assign	SYNTHESIZED_WIRE_74 = l_input[4] ~^ SYNTHESIZED_WIRE_66;

assign	SYNTHESIZED_WIRE_75 = l_input[3] ~^ SYNTHESIZED_WIRE_91;

assign	SYNTHESIZED_WIRE_76 = l_input[2] ~^ SYNTHESIZED_WIRE_68;

assign	SYNTHESIZED_WIRE_77 = l_input[1] ~^ SYNTHESIZED_WIRE_69;

assign	SYNTHESIZED_WIRE_78 = l_input[0] ~^ SYNTHESIZED_WIRE_70;

assign	SYNTHESIZED_WIRE_80 = SYNTHESIZED_WIRE_71 & SYNTHESIZED_WIRE_72 & SYNTHESIZED_WIRE_73 & SYNTHESIZED_WIRE_74;

assign	SYNTHESIZED_WIRE_81 = SYNTHESIZED_WIRE_75 & SYNTHESIZED_WIRE_76 & SYNTHESIZED_WIRE_77 & SYNTHESIZED_WIRE_78;

assign	SYNTHESIZED_WIRE_5 = l_input[5] ~^ SYNTHESIZED_WIRE_79;

assign	is_SHW = SYNTHESIZED_WIRE_80 & SYNTHESIZED_WIRE_81;

assign	SYNTHESIZED_WIRE_63 =  ~SYNTHESIZED_WIRE_91;

assign	SYNTHESIZED_WIRE_65 =  ~SYNTHESIZED_WIRE_91;

assign	SYNTHESIZED_WIRE_66 =  ~SYNTHESIZED_WIRE_91;

assign	SYNTHESIZED_WIRE_68 =  ~SYNTHESIZED_WIRE_91;

assign	SYNTHESIZED_WIRE_69 =  ~SYNTHESIZED_WIRE_91;

assign	SYNTHESIZED_WIRE_70 =  ~SYNTHESIZED_WIRE_91;

assign	SYNTHESIZED_WIRE_6 = l_input[4] ~^ SYNTHESIZED_WIRE_88;

assign	SYNTHESIZED_WIRE_7 = l_input[3] ~^ SYNTHESIZED_WIRE_89;

assign	SYNTHESIZED_WIRE_8 = l_input[2] ~^ SYNTHESIZED_WIRE_91;

assign	l_input = ASCII_Input;

endmodule
